LIBRARY ieee ;
USE ieee.std_logic_1164.all ;

ENTITY sraiBlock IS
generic(N:integer);
PORT (DATA_IN: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0) ;
	 SHIFT: IN STD_LOGIC_VECTOR(4 downto 0);
DATA_OUT: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0) ) ;
END sraiBlock ;

ARCHITECTURE Behavior OF sraiBlock IS

signal sh0, sh1, sh2, sh3, sh4, sh5, sh6, sh7, sh8, sh9, sh10, sh11, sh12, sh13, sh14, sh15, sh16, sh17, sh18, sh19, sh20, sh21, sh22,
	 sh23, sh24, sh25, sh26, sh27, sh28, sh29, sh30, sh31: STD_LOGIC_VECTOR(31 DOWNTO 0) ;
	 
	 
component mux32to1 IS
PORT (X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, X16,
	 X17, X18, X19, X20, X21, X22, X23, X24, X25, X26, X27, X28, X29, X30, X31, X32: IN STD_LOGIC_VECTOR(31 DOWNTO 0) ;
	 Sel: IN STD_LOGIC_VECTOR(4 downto 0);
Y: OUT STD_LOGIC_VECTOR(31 DOWNTO 0) ) ;
END component;

begin
sh0<=DATA_IN;
sh1<=DATA_IN(31)& DATA_IN(31 downto 1);
sh2<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31 downto 2);
sh3<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 3);
sh4<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 4);
sh5<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 5);
sh6<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 6);
sh7<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 7);
sh8<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 8);
sh9<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 9);
sh10<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 10);
sh11<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 11);
sh12<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 12);
sh13<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 13);
sh14<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 14);
sh15<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 15);
sh16<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 16);
sh17<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 17);
sh18<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 18);
sh19<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 19);
sh20<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 20);
sh21<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 21);
sh22<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 22);
sh23<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 23);
sh24<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 24);
sh25<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 25);
sh26<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 26);
sh27<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 27);
sh28<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 28);
sh29<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 29);
sh30<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31 downto 30);
sh31<=DATA_IN(31)& DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31) & DATA_IN(31);


sraimux: mux32to1 port map(sh0, sh1, sh2, sh3, sh4, sh5, sh6, sh7, sh8, sh9, sh10, sh11, sh12, sh13, sh14, sh15, sh16, sh17, sh18, sh19, sh20, sh21, sh22,
	 sh23, sh24, sh25, sh26, sh27, sh28, sh29, sh30, sh31, SHIFT, DATA_OUT);

END ARCHITECTURE;





