library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


ENTITY MUX8_1 IS
generic(N: integer);
PORT(A,B,C,D,E,F,G,H:IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
SEL:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
DOUT:OUT STD_LOGIC_VECTOR(N-1 downto 0));
END MUX8_1;

ARCHITECTURE BEH123 OF MUX8_1 IS
BEGIN
PROCESS(a,b,c,d,e,f,g,h,SEL)
BEGIN
CASE SEL IS
WHEN"000"=>DOUT<=A;
WHEN"001"=>DOUT<=B;
WHEN"010"=>DOUT<=C;
WHEN"011"=>DOUT<=D;
WHEN"100"=>DOUT<=E;
WHEN"101"=>DOUT<=F;
WHEN"110"=>DOUT<=G;
WHEN"111"=>DOUT<=H;
WHEN OTHERS=>
DOUT<=A;
END CASE;
END PROCESS;
END BEH123; 