// File ./Stage3/ALUBlock/sraiBlock.vhd translated with vhd2vl v3.0 VHDL to Verilog RTL translator
// vhd2vl settings:
//  * Verilog Module Declaration Style: 2001

// vhd2vl is Free (libre) Software:
//   Copyright (C) 2001 Vincenzo Liguori - Ocean Logic Pty Ltd
//     http://www.ocean-logic.com
//   Modifications Copyright (C) 2006 Mark Gonzales - PMC Sierra Inc
//   Modifications (C) 2010 Shankar Giri
//   Modifications Copyright (C) 2002-2017 Larry Doolittle
//     http://doolittle.icarus.com/~larry/vhd2vl/
//   Modifications (C) 2017 Rodrigo A. Melo
//
//   vhd2vl comes with ABSOLUTELY NO WARRANTY.  Always check the resulting
//   Verilog for correctness, ideally with a formal verification tool.
//
//   You are welcome to redistribute vhd2vl under certain conditions.
//   See the license (GPLv2) file included with the source for details.

// The result of translation follows.  Its copyright status should be
// considered unchanged from the original VHDL.

// no timescale needed

module sraiBlock(
input wire [N - 1:0] DATA_IN,
input wire [4:0] SHIFT,
output wire [N - 1:0] DATA_OUT
);

parameter [31:0] N = 32;



wire [31:0] sh0; wire [31:0] sh1; wire [31:0] sh2; wire [31:0] sh3; wire [31:0] sh4; wire [31:0] sh5; wire [31:0] sh6; wire [31:0] sh7; wire [31:0] sh8; wire [31:0] sh9; wire [31:0] sh10; wire [31:0] sh11; wire [31:0] sh12; wire [31:0] sh13; wire [31:0] sh14; wire [31:0] sh15; wire [31:0] sh16; wire [31:0] sh17; wire [31:0] sh18; wire [31:0] sh19; wire [31:0] sh20; wire [31:0] sh21; wire [31:0] sh22; wire [31:0] sh23; wire [31:0] sh24; wire [31:0] sh25; wire [31:0] sh26; wire [31:0] sh27; wire [31:0] sh28; wire [31:0] sh29; wire [31:0] sh30; wire [31:0] sh31;

  assign sh0 = DATA_IN;
  assign sh1 = {DATA_IN[31],DATA_IN[31:1]};
  assign sh2 = {DATA_IN[31],DATA_IN[31],DATA_IN[31:2]};
  assign sh3 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:3]};
  assign sh4 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:4]};
  assign sh5 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:5]};
  assign sh6 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:6]};
  assign sh7 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:7]};
  assign sh8 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:8]};
  assign sh9 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:9]};
  assign sh10 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:10]};
  assign sh11 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:11]};
  assign sh12 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:12]};
  assign sh13 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:13]};
  assign sh14 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:14]};
  assign sh15 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:15]};
  assign sh16 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:16]};
  assign sh17 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:17]};
  assign sh18 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:18]};
  assign sh19 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:19]};
  assign sh20 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:20]};
  assign sh21 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:21]};
  assign sh22 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:22]};
  assign sh23 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:23]};
  assign sh24 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:24]};
  assign sh25 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:25]};
  assign sh26 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:26]};
  assign sh27 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:27]};
  assign sh28 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:28]};
  assign sh29 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:29]};
  assign sh30 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31:30]};
  assign sh31 = {DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31],DATA_IN[31]};
  mux32to1 sraimux(
      sh0,
    sh1,
    sh2,
    sh3,
    sh4,
    sh5,
    sh6,
    sh7,
    sh8,
    sh9,
    sh10,
    sh11,
    sh12,
    sh13,
    sh14,
    sh15,
    sh16,
    sh17,
    sh18,
    sh19,
    sh20,
    sh21,
    sh22,
    sh23,
    sh24,
    sh25,
    sh26,
    sh27,
    sh28,
    sh29,
    sh30,
    sh31,
    SHIFT,
    DATA_OUT);


endmodule
